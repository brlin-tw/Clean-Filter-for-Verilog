`ifndef FOO
module demo();

endmodule
`endif
